module ControllerLCD(
	dataa, // operand A <always required>
	datab, // operand B <optional>
	result // result <always required>
);
	input [31:0]dataa;
	input [31:0]datab;
	output[31:0]result;
// Port Declaration
// Wire Declaration
// Integer Declaration
// Concurrent Assignment
endmodule