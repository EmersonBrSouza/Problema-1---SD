
module Main (
	clk_clk,
	push_buttons_external_connection_export,
	controllerlcd_0_conduit_end_readdata);	

	input		clk_clk;
	input	[3:0]	push_buttons_external_connection_export;
	output	[12:0]	controllerlcd_0_conduit_end_readdata;
endmodule
